module ALU
    import DEF::*;  // import package DEF in module header
(
    input alu_control_packet_t alu_control,
    input dw operand_1,
    input dw operand_2,
    output dw alu_out
);
//TODO
endmodule : ALU
