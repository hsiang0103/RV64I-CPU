module Reg_M
    import DEF::*;
(
    input logic clk,
    input logic rst,
    input dw alu_out_E,
    input dw rs2_data_E,
    input dw current_pc_E,
    output dw current_pc_M,
    output dw alu_out_M,
    output dw rs2_data_M
);
//TODO
endmodule