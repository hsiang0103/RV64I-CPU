module PC
    import DEF::*;
(
    input logic clk,
    input logic rst,
    input dw next_pc,
    input logic stall,
    output dw current_pc
);
//TODO
endmodule : PC
