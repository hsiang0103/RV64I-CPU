module Reg_E
    import DEF::*;
(
    input logic clk,
    input logic rst,
    input dw current_pc_D,
    input dw rs1_data_D,
    input dw rs2_data_D,
    input dw sext_imm_D,
    input logic stall,
    input logic jb,
    output dw current_pc_E,
    output dw rs1_data_E,
    output dw rs2_data_E,
    output dw sext_imm_E
);
//TODO
endmodule