module Reg_W
    import DEF::*;
(
    input logic clk,
    input logic rst,
    input dw alu_out_M,
    input dw ld_data_M,
    input dw current_pc_M,
    output dw current_pc_W,
    output dw alu_out_W,
    output dw ld_data_W
);
//TODO
endmodule